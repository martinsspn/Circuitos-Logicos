ENTITY pc IS
PORT()
END pc;

ARCHITECTURE arch OF pc IS
BEGIN
END arch;