ENTITY po IS
PORT()
END po;

ARCHITECTURE arch OF po IS


BEGIN

END arch;